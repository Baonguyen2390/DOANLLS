library verilog;
use verilog.vl_types.all;
entity MUL32BIT_vlg_vec_tst is
end MUL32BIT_vlg_vec_tst;
